module karatsuba64 ( input  logic        clk, input  logic        rst, input  logic        start, input  logic [63:0] A, input  logic [63:0] B, output logic [127:0] P, output logic        valid_out ); // Split 64-bit inputs logic [33:0] A_hi, A_lo, B_hi, B_lo; logic [31:0] A_hi32, A_lo32; assign A_hi32 = A >> 32; assign A_lo32 = A & 32'hFFFFFFFF; assign A_hi = {2'b0, A_hi32}; assign A_lo = {2'b0, A_lo32}; logic [31:0] B_hi32, B_lo32; assign B_hi32 = B >> 32; assign B_lo32 = B & 32'hFFFFFFFF; assign B_hi = {2'b0, B_hi32}; assign B_lo = {2'b0, B_lo32}; // Outputs of 32x32 Karatsuba units logic [67:0] z0, z1, z2; logic v0, v1, v2; logic [135:0] mid_ext, z1_ext; // extended width to prevent overflow assign mid_ext = (z2 - z1 - z0) << 32; assign z1_ext  = z1 << 64; logic [33:0] sumA, sumB; // 34-bit sum assign sumA =  A_hi + A_lo; assign sumB = B_hi + B_lo;; logic start_z0, start_z1, start_z2; // Instantiate three karatsuba34 units karatsuba34 k0 (.clk(clk), .rst(rst), .start(start_z0), .A(A_lo), .B(B_lo), .P(z0), .valid_out(v0)); karatsuba34 k1 (.clk(clk), .rst(rst), .start(start_z1), .A(A_hi), .B(B_hi), .P(z1), .valid_out(v1)); karatsuba34 k2 (.clk(clk), .rst(rst), .start(start_z2), .A(sumA), .B(sumB), .P(z2), .valid_out(v2)); // FSM states typedef enum logic [2:0] { IDLE, START_P0, WAIT_P0, START_P1, WAIT_P1, START_P2, WAIT_P2, COMBINE } state_t; state_t state; logic [127:0] P_reg; assign P = P_reg[127:0]; logic valid_reg; assign valid_out = valid_reg; always_ff @(posedge clk or posedge rst) begin if (rst) begin state <= IDLE; P_reg <= 0; valid_reg <= 0; start_z0 <= 0; start_z1 <= 0; start_z2 <= 0; end else begin // defaults start_z0 <= 0; start_z1 <= 0; start_z2 <= 0; valid_reg <= 0; case(state) IDLE: if (start) begin $display("[%0t] IDLE -> START_P0, A=%h, B=%h", $time, A, B); state <= START_P0; end // Stage 0: compute z0 = A_lo*B_lo START_P0: begin start_z0 <= 1; $display("[%0t] START_P0: A_lo=%h, B_lo=%h", $time, A_lo, B_lo); state <= WAIT_P0; end WAIT_P0: if (v0) begin $display("[%0t] WAIT_P0 done: z0=%h", $time, z0); state <= START_P1; end // Stage 1: compute z1 = A_hi*B_hi START_P1: begin start_z1 <= 1; $display("[%0t] START_P1: A_hi=%h, B_hi=%h", $time, A_hi, B_hi); state <= WAIT_P1; end WAIT_P1: if (v1) begin $display("[%0t] WAIT_P1 done: z1=%h", $time, z1); state <= START_P2; end // Stage 2: compute z2 = (A_hi+A_lo)*(B_hi+B_lo) START_P2: begin start_z2 <= 1; $display("[%0t] START_P2: sumA=%h, sumB=%h", $time, sumA, sumB); state <= WAIT_P2; end WAIT_P2: if (v2) begin $display("[%0t] WAIT_P2 done: z2=%h", $time, z2); state <= COMBINE; end // Combine results COMBINE: begin $display("[%0t] COMBINE: z0=%h, z1=%h, z2=%h", $time, z0, z1, z2); $display("[%0t] mid_ext=%h, z1_ext=%h", $time, mid_ext, z1_ext); P_reg  <= z1_ext + mid_ext + z0; // combine valid_reg <= 1; $display("[%0t] P=%h", $time, P_reg); state <= IDLE; end endcase end end endmodule